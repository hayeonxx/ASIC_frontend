module not_gate(
	input a,
	output o
);

	assign o = ~a;
endmodule
