module IOPOWER(VDD, VSS);
inout VDD;
inout VSS;

IOVDD_NS IOVDD_L1 ();
IOVDD_NS IOVDD_B1 ();
IOVDD_NS IOVDD_R1 ();
IOVDD_NS IOVDD_T1 ();

IOVSS_NS IOVSS_L1 ();
IOVSS_NS IOVSS_B1 ();
IOVSS_NS IOVSS_R1 ();
IOVSS_NS IOVSS_T1 ();

VDD_NS VDD_L1 ();
VDD_NS VDD_L2 ();
VDD_NS VDD_B1 ();
VDD_NS VDD_B2 ();
VDD_NS VDD_R1 ();
VDD_NS VDD_R2 ();
VDD_NS VDD_T1 ();
VDD_NS VDD_T2 ();

VSS_NS VSS_L1 ();
VSS_NS VSS_L2 ();
VSS_NS VSS_B1 ();
VSS_NS VSS_B2 ();
VSS_NS VSS_R1 ();
VSS_NS VSS_R2 ();
VSS_NS VSS_T1 ();
VSS_NS VSS_T2 ();

AVDD_NS AVDD_PLL1 ();
AVSS_NS AVSS_PLL1 ();
VDD_NS DVDD_PLL1 ();

AVDD_NS AVDD_PLL2 ();
AVSS_NS AVSS_PLL2 ();
VDD_NS DVDD_PLL2 ();

endmodule
